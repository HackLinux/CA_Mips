library verilog;
use verilog.vl_types.all;
entity testHW6 is
end testHW6;
